
/*
	Based on bright, hcount, vcount, turn on the bits
	Figures out the position and the color of the pixel
	Draws the pixel
*/
module bitGen ();




endmodule
