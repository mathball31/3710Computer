

/*
	Generate timing pulses at the right time
	Hsync, vsync, bright, hcount, vcount
	All about timing
	Doesn't draw anything
	
	640 x 480 pixel screen
*/
module VGAControl ();



endmodule
